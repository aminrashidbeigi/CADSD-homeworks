----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 10/31/2017 11:33:03 AM
-- Design Name: 
-- Module Name: counter - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
--use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity counter is
    port(
    clk, rst: in std_logic;
    module: in integer := 4;
    output: out std_logic_vector(5 downto 0)
    );
end counter;

architecture Behavioral of counter is

component counter_mod_m is
    generic(
    module: std_logic_vector(5 downto 0)
    );
    port(
    clk, rst: in std_logic;
    output: out std_logic_vector(5 downto 0)
    );
end component;


begin
    counter_module: counter_mod_m generic map (std_logic_vector(to_unsigned(module, 6))) port map (clk,rst,output);
    
end Behavioral;
